`timescale 1ns/1ns
`include "../processador/mpc.v"


module mpc_tb;
    reg [15:0]pcp; 
    reg [15:0]pcj; 
    reg choice;
    wire[15:0] out;

    mpc mux( 
        pcp,
        pcj,
        choice,
        out
    );

    initial begin
        $monitor("PCp = %d, PCJ = %d, choice = %b, out = %d", pcp, pcj, choice, out);
        //$dumpfile ("testbench/ACControl.vcd");    
	    //$dumpvars(0, ACControl_tb);

        pcp = 16'b0000000000000010;
        pcj = 16'b0000000001111100;
        choice = 1;

        #20
        pcp = 16'b0000000000001110;
        pcj = 16'b0000000001111100;
        choice = 0;


        #20
        $monitor("test completed");
    end

endmodule